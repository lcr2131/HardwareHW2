testbench yo