top file, real big