//Author: Leonard Robinson
class;


	function void golden_result;
	  $display();
	end function

	function bit check_result();
		return;
	end function
end class

program (iffc.bench x) //iffc is the interface of the flip flop class

	initial begin
	 repeat
	  $display
	  $display
	 end //end repeat
	end //end initial
	

end program