module cam_module(ifc.dut_cam  d)
  


  endmodule 

