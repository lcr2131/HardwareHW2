//Author: Leonard Robinson